
module dual_port_ram #(parameter ADDR_WIDTH = 6,parameter DATA_WIDTH = 16,parameter DEPTH = 64)   
  							(input [DATA_WIDTH :0] data_a, data_b,
                         	 input [ADDR_WIDTH-1:0] addr_a, addr_b,
                        	 input we_a, we_b, clk,
                             output reg [DATA_WIDTH-1:0] q_a, q_b );

 reg [DATA_WIDTH:0] ram[DEPTH:0];
	
// Port A
always @ (posedge clk)
    begin
      if (we_a) 
        begin
          ram[addr_a] <= data_a;
          q_a <= data_a;
        end
      else 
        q_a <= ram[addr_a];        
    end
	
// Port B
always @ (posedge clk)
	begin
		if (we_b)
          begin
              ram[addr_b] <= data_b;
              q_b <= data_b;
          end
		else
              q_b <= ram[addr_b];
	end
  
endmodule
